module Issue_2_2 (
    input clk_50MHz_i,
    input clk_100MHz_i,
    input idat
);

endmodule